module pll_m1t(
    input areset,
    output inclk0,
    output c0,
    output locked
);

    // Just a black box

endmodule : pll_m1t