module Toplevel_m1t #(
    IS_TESTBENCH = 0
)(
    input  wire        clk,
    input  wire        async_rst,
    //input  wire [15:0] gpi,
    //output wire [15:0] gpo
    output wire [7:0] gpo
);

    wire [15:0] gpi = 'h0;

    wire gen_clk;
    generate
        if(IS_TESTBENCH) begin
            assign gen_clk = clk;
        end else begin
            pll_m1t pll (
            .areset(!async_rst),
            .inclk0(clk),
            .c0(gen_clk),
            .locked()
            );
        end
    endgenerate
    

    reg [15:0] irom [2047:0];
    reg [15:0] irom_buffer;

    initial begin
        if(IS_TESTBENCH) $readmemh("/mnt/e/programacion/systemverilog/MINT/M1/rtl/test_programs/test.txt", irom);
		else $readmemh("E:/programacion/systemverilog/MINT/M1/rtl/test_programs/test.txt", irom);
    end

    always_ff @(posedge clk) begin
        if(rom_req) begin
            irom_buffer <= irom[inst_addr[10:0]];
        end
    end

    always_ff @(posedge clk) begin
        rst_buffer0 <= !async_rst;
        rst_buffer1 <= rst_buffer0;
    end

    reg rst_buffer0 = 'b1;
    reg rst_buffer1 = 'b1;
    wire sync_rst = rst_buffer0 && rst_buffer1;

    wire rom_req;
    wire [14:0] inst_addr;

    wire [14:0] mem_address_out;
    wire [1:0]  mem_mask_out;
    wire [1:0]  mem_read_fnc_type;
    wire [15:0] mem_data_out;
    wire [1:0]  mem_mode;
    wire        mem_enable;
    wire [3:0]  mem_wb_dest;
    wire        mem_input_ready;
    wire [15:0] mem_data_in;
    wire [3:0]  mem_wb_dest_in;
    wire        mem_read_ack;
    wire        mem_available;
    wire        mem_idle;

    Core_m1 Core (
        .clk                (gen_clk),
        .clk_en             ('b1),
        .sync_rst           (sync_rst),
        .icache_miss        ('b0),
        .instruction_in     (irom_buffer),
        .icache_req         (rom_req),
        .inst_address_out   (inst_addr),
        .mem_address_out    (mem_address_out),
        .mem_mask_out       (mem_mask_out),
        .mem_read_fnc_type  (mem_read_fnc_type),
        .mem_data_out       (mem_data_out),
        .mem_mode           (mem_mode),
        .mem_enable         (mem_enable),
        .mem_wb_dest        (mem_wb_dest),
        .mem_input_ready    (mem_input_ready),
        .mem_data_in        (mem_data_in),
        .mem_wb_dest_in     (mem_wb_dest_in),
        .mem_read_ack       (mem_read_ack),
        .mem_available      (mem_available),
        .mem_idle           (mem_idle)
    );

    MemoryController_m1t MemoryController (
        .clk                        (gen_clk),
        .clk_en                     ('b1),
        .sync_rst                   (sync_rst),
        .core_mem_address_out       (mem_address_out),
        .core_mem_mask_out          (mem_mask_out),
        .core_mem_read_fnc_type     (mem_read_fnc_type),
        .core_mem_data_out          (mem_data_out),
        .core_mem_mode              (mem_mode),
        .core_mem_enable            (mem_enable && !mem_mode[1]),
        .core_mem_wb_dest           (mem_wb_dest),
        .core_mem_input_ready       (mem_input_ready),
        .core_mem_data_in           (mem_data_in),
        .core_mem_wb_dest_in        (mem_wb_dest_in),
        .core_mem_read_ack          (mem_read_ack),
        .core_mem_available         (mem_available),
        .core_mem_idle              (mem_idle),
        .gpo_bank                   (gpo),
        .gpi_bank                   (gpi)
    );

endmodule : Toplevel_m1t